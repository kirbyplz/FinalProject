module snn_core(addr_input_unit, digit, done, start, q_input);

input start, q_input;
output done;
output [3:0] digit;
output [9:0] addr_input_unit;




endmodule
